`include "Lab4.v"

module TestBench();

  initial
  begin
    #10

    $finish
  end

endmodule
