module Lab3();
endmodule
